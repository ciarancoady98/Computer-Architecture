---------------------------------------------------------------------------------- 
-- Engineer: Ciaran Coady
-- Module Name: Full_Adder_tb
-- Project Name: Computer Architecture
----------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

ENTITY Full_Adder_tb IS
END Full_Adder_tb;
 
ARCHITECTURE behavior OF Full_Adder_tb is
 
    -- Component Declaration for the Unit Under Test (UUT)
    component Full_Adder
    Port ( In1 : in STD_LOGIC;
           In2 : in STD_LOGIC;
           C_in : in STD_LOGIC;
           Sum : out STD_LOGIC;
           C_out : out STD_LOGIC);
    end component;
    

   --Inputs
   signal In1_signal : STD_LOGIC;
   signal In2_signal : STD_LOGIC;
   signal C_in_signal : STD_LOGIC;

 	--Outputs
   signal Sum_signal : STD_LOGIC;
   signal C_out_signal : STD_LOGIC;
   
   --Clock
   constant Clk_period : time := 40 ns;
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: Full_Adder PORT MAP (
          In1 => In1_signal,
          In2 => In2_signal,
          C_in => C_in_signal,
          Sum => Sum_signal,
          C_out => C_out_signal
        );

   stim_proc: process
   begin	
        
      wait for Clk_period;
      --Cin = 0, 0+0=0, Cout = 0
      In1_signal <= '0';
      In2_signal <= '0';
      C_in_signal <= '0';
      
      wait for Clk_period;
      
      --Cin = 0, 1+0=1, Cout = 0
      In1_signal <= '1';
      In2_signal <= '0';
      C_in_signal <= '0';
      
      wait for Clk_period;	
      
      --Cin = 0, 1+1=0, Cout = 1
      In1_signal <= '1';
      In2_signal <= '1';
      C_in_signal <= '0';
      
      wait for Clk_period;
      	
      --Cin = 1, 0+0=1, Cout = 0
      In1_signal <= '0';
      In2_signal <= '0';
      C_in_signal <= '1';
      
      wait for Clk_period;	
      
      --Cin = 1, 0+1=0, Cout = 1
      In1_signal <= '0';
      In2_signal <= '1';
      C_in_signal <= '1';
      
      wait for Clk_period;
      
      --Cin = 1, 1+1=1, Cout = 1
      In1_signal <= '1';
      In2_signal <= '1';
      C_in_signal <= '1';
     
      wait for Clk_period;
     
   end process;

END;