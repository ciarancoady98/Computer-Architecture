---------------------------------------------------------------------------------- 
-- Engineer: Ciaran Coady
-- Module Name: Ripple_Adder_16bit_tb
-- Project Name: Computer Architecture
----------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

ENTITY Ripple_Adder_16bit_tb IS
END Ripple_Adder_16bit_tb;
 
ARCHITECTURE behavior OF Ripple_Adder_16bit_tb is
 
    -- Component Declaration for the Unit Under Test (UUT)
    component Ripple_Adder_16bit
    Port ( X : in STD_LOGIC_VECTOR (15 downto 0);
           Y : in STD_LOGIC_VECTOR (15 downto 0);
           C_in : in STD_LOGIC;
           Z : out STD_LOGIC_VECTOR (15 downto 0);
           C_out : out STD_LOGIC);
    end component;
    

   --Inputs
   signal X_signal : STD_LOGIC_VECTOR (15 downto 0);
   signal Y_signal : STD_LOGIC_VECTOR (15 downto 0);
   signal C_in_signal : STD_LOGIC;

 	--Outputs
   signal Z_signal : STD_LOGIC_VECTOR (15 downto 0);
   signal C_out_signal : STD_LOGIC;
   
   --Clock
   constant Clk_period : time := 40 ns;
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: Ripple_Adder_16bit PORT MAP (
          X => X_signal,
          Y => Y_signal,
          C_in => C_in_signal,
          Z => Z_signal,
          C_out => C_out_signal
        );

   stim_proc: process
   begin	
        
      wait for Clk_period*3;
      
      --Cin = 0, 0+0=0, Cout = 0
      X_signal <= "0000000000000000";
      Y_signal <= "0000000000000000";
      C_in_signal <= '0';
      
      wait for Clk_period*3;
      
      --Cin = 0, 1+0=1, Cout = 0
      X_signal <= "0000000000000001";
      
      wait for Clk_period*3;	
      
      --Cin = 0, 1+1=2, Cout = 0
      X_signal <= "0000000000000001";
      Y_signal <= "0000000000000001";
      
      wait for Clk_period*3;
      	
      --Cin = 1, 1+1=3, Cout = 0
      C_in_signal <= '1';
      
      wait for Clk_period*3;
      
      C_in_signal <= '0';
      
      wait for Clk_period*3;
      
      --Cin = 1, FFFE+FFFF=0, Cout = 1
      C_in_signal <= '0';
      X_signal <= "1111111111111110";
      Y_signal <= "1111111111111111";
     
      wait for Clk_period*3;
     
   end process;

END;