---------------------------------------------------------------------------------- 
-- Engineer: Ciaran Coady
-- Module Name: Memory_512
-- Project Name: Computer Architecture
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity Memory_512 is
    Port ( Address_in : in STD_LOGIC_VECTOR (15 downto 0);
           Data_in : in  STD_LOGIC_VECTOR (15 downto 0);
           Clk : in STD_LOGIC;
           MW : in  STD_LOGIC;
           Data_out : out  STD_LOGIC_VECTOR (15 downto 0));
end Memory_512;

architecture Behavioral of Memory_512 is

type mem_array is array(0 to 511) of std_logic_vector(15 downto 0);

begin

mem_process: process (Address_in, Data_in,Clk)

variable data_mem : mem_array := (

--			               		          Instructions					Instruction Code			
--																        Opcode  DR  SA  SB

"0000000010010011", 					--ADI R2, R2, #3				0000000 010 010 011 		
"0000101011010010", 					--ADD R3, R2, R2  				0000101 011 010 010 		
"0000000001001010", 					--ADI R1, R1, #2				0000000 001 001 010		    
"0000001111010000", 					--LD  R7, Memory[R2]			0000001 111 010 000
"0000101011011011", 					--ADD R3, R3, R3				0000101 011 011 011		    	    
"0000100011011000", 					--NOT R3, R3      			    0000100 011 011 000	
"0000111100100100", 					--SR  R4, R4, R4		    	0000111 100 100 100			    

X"0000", X"0000", X"0000",X"0000",
X"0000", X"0000", X"0000",X"0000",
X"0000",

X"0000", X"0000", X"0000",X"0000",		
X"0000", X"0000", X"0000",X"0000",
X"0000", X"0000", X"0000",X"0000",
X"0000", X"0000", X"0000",X"0000",

X"0000", X"0000", X"0000",X"0000",		
X"0000", X"0000", X"0000",X"0000",
X"0000", X"0000", X"0000",X"0000",
X"0000", X"0000", X"0000",X"0000",

X"0000", X"0000", X"0000",X"0000",		
X"0000", X"0000", X"0000",X"0000",
 X"0000", X"0000",X"0000",X"0000",
X"0000", X"0000", X"0000",X"0000",

X"0000", X"0000", X"0000",X"0000",		
X"0000", X"0000", X"0000",X"0000",
 X"0000", X"0000",X"0000",X"0000",
X"0000", X"0000", X"0000",X"0000",

X"0000", X"0000", X"0000",X"0000",		
X"0000", X"0000", X"0000",X"0000",
 X"0000", X"0000",X"0000",X"0000",
X"0000", X"0000", X"0000",X"0000",

X"0000", X"0000", X"0000",X"0000",	
X"0000", X"0000", X"0000",X"0000",
 X"0000", X"0000",X"0000",X"0000",
X"0000", X"0000", X"0000",X"0000",

X"0000", X"0000", X"0000",X"0000",	
X"0000", X"0000", X"0000",X"0000",
 X"0000", X"0000",X"0000",X"0000",
X"0000", X"0000", X"0000",X"0000",

X"0000", X"0000", X"0000",X"0000",		
X"0000", X"0000", X"0000",X"0000",
 X"0000", X"0000",X"0000",X"0000",
X"0000", X"0000", X"0000",X"0000",

X"0000", X"0000", X"0000",X"0000",		
X"0000", X"0000", X"0000",X"0000",
 X"0000", X"0000",X"0000",X"0000",
X"0000", X"0000", X"0000",X"0000",

X"0000", X"0000", X"0000",X"0000",	
X"0000", X"0000", X"0000",X"0000",
 X"0000", X"0000",X"0000",X"0000",
X"0000", X"0000", X"0000",X"0000",

X"0000", X"0000", X"0000",X"0000",
X"0000", X"0000", X"0000",X"0000",
 X"0000", X"0000",X"0000",X"0000",
X"0000", X"0000", X"0000",X"0000",

X"0000", X"0000", X"0000",X"0000",	
X"0000", X"0000", X"0000",X"0000",
 X"0000", X"0000",X"0000",X"0000",
X"0000", X"0000", X"0000",X"0000",

X"0000", X"0000", X"0000",X"0000",	
X"0000", X"0000", X"0000",X"0000",
 X"0000", X"0000",X"0000",X"0000",
X"0000", X"0000", X"0000",X"0000",

X"0000", X"0000", X"0000",X"0000",	
X"0000", X"0000", X"0000",X"0000",
 X"0000", X"0000",X"0000",X"0000",
X"0000", X"0000", X"0000",X"0000",

X"0000", X"0000", X"0000",X"0000",	
X"0000", X"0000", X"0000",X"0000",
 X"0000", X"0000",X"0000",X"0000",
X"0000", X"0000", X"0000",X"0000",

X"0000", X"0000", X"0000",X"0000",	
X"0000", X"0000", X"0000",X"0000",
 X"0000", X"0000",X"0000",X"0000",
X"0000", X"0000", X"0000",X"0000",

X"0000", X"0000", X"0000",X"0000",
X"0000", X"0000", X"0000",X"0000",
 X"0000", X"0000",X"0000",X"0000",
X"0000", X"0000", X"0000",X"0000",

X"0000", X"0000", X"0000",X"0000",
X"0000", X"0000", X"0000",X"0000",
 X"0000", X"0000",X"0000",X"0000",
X"0000", X"0000", X"0000",X"0000",

X"0000", X"0000", X"0000",X"0000",
X"0000", X"0000", X"0000",X"0000",
 X"0000", X"0000",X"0000",X"0000",
X"0000", X"0000", X"0000",X"0000",

X"0000", X"0000", X"0000",X"0000",	
X"0000", X"0000", X"0000",X"0000",
 X"0000", X"0000",X"0000",X"0000",
X"0000", X"0000", X"0000",X"0000",

X"0000", X"0000", X"0000",X"0000",	
X"0000", X"0000", X"0000",X"0000",
 X"0000", X"0000",X"0000",X"0000",
X"0000", X"0000", X"0000",X"0000",

X"0000", X"0000", X"0000",X"0000",
X"0000", X"0000", X"0000",X"0000",
 X"0000", X"0000",X"0000",X"0000",
X"0000", X"0000", X"0000",X"0000",

X"0000", X"0000", X"0000",X"0000",
X"0000", X"0000", X"0000",X"0000",
 X"0000", X"0000",X"0000",X"0000",
X"0000", X"0000", X"0000",X"0000",

X"0000", X"0000", X"0000",X"0000",
X"0000", X"0000", X"0000",X"0000",
 X"0000", X"0000",X"0000",X"0000",
X"0000", X"0000", X"0000",X"0000",

X"0000", X"0000", X"0000",X"0000",
X"0000", X"0000", X"0000",X"0000",
 X"0000", X"0000",X"0000",X"0000",
X"0000", X"0000", X"0000",X"0000",

X"0000", X"0000", X"0000",X"0000",
X"0000", X"0000", X"0000",X"0000",
 X"0000", X"0000",X"0000",X"0000",
X"0000", X"0000", X"0000",X"0000",

X"0000", X"0000", X"0000",X"0000",
X"0000", X"0000", X"0000",X"0000",
 X"0000", X"0000",X"0000",X"0000",
X"0000", X"0000", X"0000",X"0000",

X"0000", X"0000", X"0000",X"0000",
X"0000", X"0000", X"0000",X"0000",
 X"0000", X"0000",X"0000",X"0000",
X"0000", X"0000", X"0000",X"0000",

X"0000", X"0000", X"0000",X"0000",
X"0000", X"0000", X"0000",X"0000",
 X"0000", X"0000",X"0000",X"0000",
X"0000", X"0000", X"0000",X"0000",

X"0000", X"0000", X"0000",X"0000",
X"0000", X"0000", X"0000",X"0000",
 X"0000", X"0000",X"0000",X"0000",
X"0000", X"0000", X"0000",X"0000",

X"0000", X"0000", X"0000",X"0000",
X"0000", X"0000", X"0000",X"0000",
 X"0000", X"0000",X"0000",X"0000",
X"0000", X"0000", X"0000",X"0000"  );
variable addr:integer;

begin -- the following type conversion function is in std_logic_arith

addr:= to_integer(unsigned(Address_in(2 downto 0)));

if MW ='1' then
data_mem(addr) := Data_in;
elsif MW = '0' then
Data_out <= data_mem(addr) after 1 ns;
end if;
end process;

end Behavioral;
