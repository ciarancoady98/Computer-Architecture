---------------------------------------------------------------------------------- 
-- Engineer: Ciaran Coady
-- Module Name: Multiplexer_16to1
-- Project Name: Computer Architecture
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity Multiplexer_16to1 is
    Port ( S0 : in  STD_LOGIC;
           S1 : in  STD_LOGIC;
           S2 : in  STD_LOGIC;
           S3 : in  STD_LOGIC;
           In0 : in  STD_LOGIC_VECTOR (15 downto 0);
           In1 : in  STD_LOGIC_VECTOR (15 downto 0);
           In2 : in  STD_LOGIC_VECTOR (15 downto 0);
           In3 : in  STD_LOGIC_VECTOR (15 downto 0);
           In4 : in  STD_LOGIC_VECTOR (15 downto 0);
           In5 : in  STD_LOGIC_VECTOR (15 downto 0);
           In6 : in  STD_LOGIC_VECTOR (15 downto 0);
           In7 : in  STD_LOGIC_VECTOR (15 downto 0);
           In8 : in  STD_LOGIC_VECTOR (15 downto 0);
           In9 : in  STD_LOGIC_VECTOR (15 downto 0);
           In10 : in  STD_LOGIC_VECTOR (15 downto 0);
           In11 : in  STD_LOGIC_VECTOR (15 downto 0);
           In12 : in  STD_LOGIC_VECTOR (15 downto 0);
           In13 : in  STD_LOGIC_VECTOR (15 downto 0);
           In14 : in  STD_LOGIC_VECTOR (15 downto 0);
           In15 : in  STD_LOGIC_VECTOR (15 downto 0);
           Z : out STD_LOGIC_VECTOR (15 downto 0));
end Multiplexer_16to1;

architecture Behavioral of Multiplexer_16to1 is

begin

Z <= In0 after 5 ns when (S0='0' and S1='0' and S2='0' and S3='0') else
In1 after 5 ns when (S0='1' and S1='0' and S2='0' and S3='0') else
In2 after 5 ns when (S0='0' and S1='1' and S2='0' and S3='0') else
In3 after 5 ns when (S0='1' and S1='1' and S2='0' and S3='0') else
In4 after 5 ns when (S0='0' and S1='0' and S2='1' and S3='0') else
In5 after 5 ns when (S0='1' and S1='0' and S2='1' and S3='0') else
In6 after 5 ns when (S0='0' and S1='1' and S2='1' and S3='0') else
In7 after 5 ns when (S0='1' and S1='1' and S2='1' and S3='0') else
In8 after 5 ns when (S0='0' and S1='0' and S2='0' and S3='1') else
In9 after 5 ns when (S0='1' and S1='0' and S2='0' and S3='1') else
In10 after 5 ns when (S0='0' and S1='1' and S2='0' and S3='1') else
In11 after 5 ns when (S0='1' and S1='1' and S2='0' and S3='1') else
In12 after 5 ns when (S0='0' and S1='0' and S2='1' and S3='1') else
In13 after 5 ns when (S0='1' and S1='0' and S2='1' and S3='1') else
In14 after 5 ns when (S0='0' and S1='1' and S2='1' and S3='1') else
In15 after 5 ns when (S0='1' and S1='1' and S2='1' and S3='1') else
"0000000000000000" after 5 ns;

end Behavioral;
